CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
300 230 30 200 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
40 C:\Users\baris\Desktop\May�s\cm6\BOM.DAT
0 7
38 96 1498 799
177209362 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 651 196 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 S
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 642 478 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
1 R
14 -10 21 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 516 480 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 CP
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 431 372 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6153 0 0
0
0
14 Logic Display~
6 854 251 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 813 252 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
9 2-In AND~
219 525 282 0 3 22
0 4 6 5
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9914 0 0
0
0
5 4027~
219 655 415 0 7 32
0 9 4 7 4 8 6 2
0
0 0 4720 0
4 4027
7 -60 35 -52
1 B
29 -61 36 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0
65 0 0 0 2 2 1 0
1 U
3747 0 0
0
0
5 4027~
219 653 307 0 7 32
0 9 5 7 5 8 10 3
0
0 0 4720 0
4 4027
7 -60 35 -52
1 A
29 -61 36 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 219563378
65 0 0 512 2 1 1 0
1 U
3549 0 0
0
0
14
7 1 2 0 0 4224 0 8 5 0 0 3
679 379
854 379
854 269
7 1 3 0 0 8320 0 9 6 0 0 3
677 271
677 270
813 270
0 4 4 0 0 8320 0 0 8 4 0 3
461 372
461 397
631 397
0 2 4 0 0 0 0 0 8 8 0 4
459 372
557 372
557 379
631 379
4 0 5 0 0 4224 0 9 0 0 6 3
629 289
568 289
568 282
3 2 5 0 0 0 0 7 9 0 0 4
546 282
580 282
580 271
629 271
6 2 6 0 0 12416 0 8 7 0 0 6
685 397
752 397
752 194
480 194
480 291
501 291
1 1 4 0 0 0 0 4 7 0 0 4
443 372
460 372
460 273
501 273
0 3 7 0 0 8192 0 0 9 10 0 5
517 388
517 312
614 312
614 280
629 280
1 3 7 0 0 8320 0 3 8 0 0 3
517 467
517 388
631 388
0 5 8 0 0 8320 0 0 9 12 0 5
654 446
719 446
719 321
653 321
653 313
1 5 8 0 0 0 0 2 8 0 0 4
643 465
643 446
655 446
655 421
0 1 9 0 0 8320 0 0 8 14 0 5
653 229
602 229
602 335
655 335
655 358
1 1 9 0 0 0 0 1 9 0 0 3
651 208
653 208
653 250
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
