CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
1958 96 3418 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
56 C:\Users\baris\Desktop\Yeni klas�r (2)\May�s\cm6\BOM.DAT
0 7
1958 96 3418 799
143654930 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 348 205 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 S
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 351 105 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 R
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 619 368 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 619 290 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
10 2-In NAND~
219 487 387 0 3 22
0 3 4 5
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5394 0 0
0
0
10 2-In NAND~
219 471 311 0 3 22
0 2 5 4
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7734 0 0
0
0
9 2-In NOR~
219 471 197 0 3 22
0 6 2 7
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9914 0 0
0
0
9 2-In NOR~
219 468 108 0 3 22
0 3 7 6
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3747 0 0
0
0
14 Logic Display~
6 720 217 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
14 Logic Display~
6 718 125 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 Q
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7931 0 0
0
0
12
0 1 2 0 0 4224 0 0 6 11 0 3
388 205
388 302
447 302
0 1 3 0 0 4224 0 0 5 12 0 3
400 105
400 378
463 378
0 2 4 0 0 8192 0 0 5 6 0 5
528 311
528 339
412 339
412 396
463 396
0 2 5 0 0 8320 0 0 6 5 0 5
561 386
561 357
429 357
429 320
447 320
3 1 5 0 0 0 0 5 3 0 0 3
514 387
514 386
619 386
3 1 4 0 0 4224 0 6 4 0 0 3
498 311
619 311
619 308
1 0 6 0 0 12288 0 7 0 0 9 5
458 188
443 188
443 142
538 142
538 108
0 2 7 0 0 8192 0 0 8 10 0 5
552 197
552 166
424 166
424 117
455 117
3 1 6 0 0 4224 0 8 10 0 0 4
507 108
653 108
653 143
718 143
3 1 7 0 0 4224 0 7 9 0 0 4
510 197
652 197
652 235
720 235
1 2 2 0 0 128 0 1 7 0 0 4
360 205
391 205
391 206
458 206
1 1 3 0 0 128 0 2 8 0 0 4
363 105
400 105
400 99
455 99
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
