CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
60 10 30 200 9
44 104 1504 807
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
34 C:\Users\baris\Desktop\cm6\BOM.DAT
0 7
44 104 1504 807
143654930 0
0
6 Title:
5 Name:
0
0
0
9
13 Logic Switch~
5 222 242 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 Z
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 223 200 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 Y
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 227 125 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
14 Logic Display~
6 554 181 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 C
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
2 +V
167 373 262 0 1 3
0 4
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5394 0 0
0
0
7 Ground~
168 352 276 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
14 Logic Display~
6 554 133 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 S
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9914 0 0
0
0
9 Inverter~
13 328 128 0 2 22
0 5 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3747 0 0
0
0
4 4539
219 433 164 0 14 29
0 5 9 9 5 2 4 5 10 2
2 6 7 3 8
0
0 0 13040 0
4 4539
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 4 5 6 1 13 12 11 10
15 2 14 9 7 3 4 5 6 1
13 12 11 10 15 2 14 9 7 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
14
13 1 3 0 0 8320 0 9 4 0 0 3
465 191
465 199
554 199
1 6 4 0 0 8320 0 5 9 0 0 4
373 271
391 271
391 173
401 173
9 0 2 0 0 4096 0 9 0 0 8 2
401 200
352 200
7 0 5 0 0 4224 0 9 0 0 14 3
401 182
303 182
303 152
1 11 6 0 0 12416 0 2 9 0 0 4
235 200
256 200
256 218
401 218
1 12 7 0 0 4224 0 1 9 0 0 4
234 242
374 242
374 227
401 227
0 10 2 0 0 0 0 0 9 8 0 3
352 211
352 209
395 209
1 5 2 0 0 4224 0 6 9 0 0 3
352 270
352 164
395 164
14 1 8 0 0 4224 0 9 7 0 0 5
465 146
528 146
528 156
554 156
554 151
0 1 5 0 0 0 0 0 9 14 0 3
388 155
388 128
401 128
0 2 9 0 0 12288 0 0 9 12 0 4
362 128
376 128
376 137
401 137
2 3 9 0 0 12416 0 8 9 0 0 4
349 128
362 128
362 146
401 146
0 1 5 0 0 0 0 0 8 14 0 3
303 125
303 128
313 128
1 4 5 0 0 128 0 3 9 0 0 4
239 125
303 125
303 155
401 155
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
