CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
320 150 30 120 9
38 96 1498 799
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
40 C:\Users\baris\Desktop\May�s\cm6\BOM.DAT
0 7
38 96 1498 799
177209362 0
0
6 Title:
5 Name:
0
0
0
25
5 4011~
219 1034 607 0 3 22
0 4 5 7
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 4 0
1 U
8953 0 0
0
0
5 4011~
219 1040 549 0 3 22
0 3 2 6
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 4 0
1 U
4441 0 0
0
0
9 Inverter~
13 1127 549 0 2 22
0 6 10
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
3618 0 0
0
0
9 Inverter~
13 1125 607 0 2 22
0 7 9
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
6153 0 0
0
0
5 4011~
219 1201 575 0 3 22
0 10 9 8
0
0 0 608 0
4 4011
-7 -24 21 -16
3 U4D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 4 2 0
1 U
5394 0 0
0
0
14 Logic Display~
6 1310 554 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7734 0 0
0
0
13 Logic Switch~
5 838 352 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
9 2 23 10
2 E1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 784 351 0 1 11
0 12
0
0 0 21360 90
2 0V
11 0 25 8
2 E2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 726 352 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 E3
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 647 288 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 Z
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 644 246 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 Y
-2 -26 5 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 641 201 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
1 X
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8903 0 0
0
0
14 Logic Display~
6 1256 410 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 C1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 1286 425 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 S
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
5 4011~
219 1189 443 0 3 22
0 10 9 8
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 3 2 0
1 U
7668 0 0
0
0
9 Inverter~
13 1101 478 0 2 22
0 7 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
4718 0 0
0
0
9 Inverter~
13 1103 420 0 2 22
0 6 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
3874 0 0
0
0
5 4011~
219 1020 427 0 3 22
0 3 2 6
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 431425072
65 0 0 0 4 2 2 0
1 U
6671 0 0
0
0
5 4011~
219 1022 486 0 3 22
0 4 5 7
0
0 0 624 0
4 4011
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 280430137
65 0 0 0 4 1 2 0
1 U
3789 0 0
0
0
7 74LS138
19 901 472 0 14 29
0 16 15 14 11 12 13 3 23 24
2 25 4 5 26
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
2 U3
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
4871 0 0
0
0
14 Logic Display~
6 1105 289 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 C
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 512 0 0 0 0
1 L
3750 0 0
0
0
10 4-In NAND~
219 1050 310 0 5 22
0 28 29 30 31 32
0
0 0 624 0
6 74LS20
-21 -28 21 -20
3 U2B
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 515311159
65 0 0 512 2 2 1 0
1 U
8778 0 0
0
0
10 4-In NAND~
219 1050 242 0 5 22
0 18 19 20 21 17
0
0 0 624 0
6 74LS20
-21 -28 21 -20
3 U2A
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 515311159
65 0 0 0 2 1 1 0
1 U
538 0 0
0
0
14 Logic Display~
6 1086 203 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 S
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6843 0 0
0
0
7 74LS138
19 931 249 0 14 29
0 16 15 14 11 12 13 18 33 34
19 35 20 21 36
0
0 0 5104 0
7 74LS138
-25 -61 24 -53
2 U1
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 512 1 0 0 0
1 U
3136 0 0
0
0
40
11 2 0 0 0 0 0 20 1 0 0 4
939 481
963 481
963 616
1010 616
9 1 0 0 0 0 0 20 1 0 0 4
939 463
957 463
957 598
1010 598
8 2 0 0 0 0 0 20 2 0 0 4
939 454
973 454
973 558
1016 558
0 1 0 0 0 0 0 0 2 16 0 3
980 418
980 540
1016 540
11 4 0 0 0 0 0 25 22 0 0 4
969 258
988 258
988 324
1026 324
9 3 0 0 0 0 0 25 22 0 0 4
969 240
979 240
979 315
1026 315
8 2 0 0 0 0 0 25 22 0 0 4
969 231
995 231
995 306
1026 306
0 1 0 0 0 0 0 0 22 31 0 3
1000 222
1000 297
1026 297
3 1 6 0 0 16 0 2 3 0 0 2
1067 549
1112 549
3 1 7 0 0 16 0 1 4 0 0 2
1061 607
1110 607
3 1 8 0 0 16 0 5 6 0 0 4
1228 575
1295 575
1295 572
1310 572
2 2 9 0 0 16 0 4 5 0 0 4
1146 607
1179 607
1179 584
1177 584
2 1 10 0 0 16 0 3 5 0 0 4
1148 549
1175 549
1175 566
1177 566
5 1 0 0 0 0 0 22 21 0 0 3
1077 310
1105 310
1105 307
10 2 2 0 0 8320 0 20 18 0 0 4
939 472
969 472
969 436
996 436
7 1 3 0 0 12416 0 20 18 0 0 4
939 445
965 445
965 418
996 418
12 1 4 0 0 4224 0 20 19 0 0 4
939 490
973 490
973 477
998 477
13 2 5 0 0 4224 0 20 19 0 0 4
939 499
971 499
971 495
998 495
3 1 6 0 0 12416 0 18 17 0 0 4
1047 427
1060 427
1060 420
1088 420
3 1 7 0 0 12416 0 19 16 0 0 4
1049 486
1062 486
1062 478
1086 478
3 1 8 0 0 4224 0 15 14 0 0 2
1216 443
1286 443
2 2 9 0 0 4224 0 16 15 0 0 4
1122 478
1155 478
1155 452
1165 452
2 1 10 0 0 4224 0 17 15 0 0 4
1124 420
1151 420
1151 434
1165 434
0 4 11 0 0 4224 0 0 20 39 0 3
820 267
820 490
869 490
0 5 12 0 0 4224 0 0 20 40 0 3
830 276
830 499
863 499
0 6 13 0 0 4224 0 0 20 38 0 3
852 285
852 508
863 508
0 3 14 0 0 4224 0 0 20 35 0 3
858 240
858 463
869 463
0 2 15 0 0 4224 0 0 20 36 0 3
868 231
868 454
869 454
0 1 16 0 0 4224 0 0 20 37 0 3
876 222
876 445
869 445
5 1 17 0 0 8320 0 23 24 0 0 3
1077 242
1086 242
1086 221
7 1 18 0 0 4224 0 25 23 0 0 4
969 222
1015 222
1015 229
1026 229
10 2 19 0 0 12416 0 25 23 0 0 4
969 249
985 249
985 238
1026 238
12 3 20 0 0 4224 0 25 23 0 0 4
969 267
998 267
998 247
1026 247
13 4 21 0 0 4224 0 25 23 0 0 4
969 276
1006 276
1006 256
1026 256
1 3 14 0 0 128 0 10 25 0 0 6
659 288
708 288
708 260
770 260
770 240
899 240
1 2 15 0 0 128 0 11 25 0 0 4
656 246
722 246
722 231
899 231
1 1 16 0 0 128 0 12 25 0 0 4
653 201
828 201
828 222
899 222
1 6 13 0 0 128 0 7 25 0 0 3
839 339
839 285
893 285
1 4 11 0 0 128 0 9 25 0 0 3
727 339
727 267
899 267
1 5 12 0 0 128 0 8 25 0 0 3
785 338
785 276
893 276
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
